module s344 (.Z(GND,VDD,CLK,A0,A1,A2,A3,B0,B1,B2,B3,CNTVCO2,CNTVCON2,P0,P1,P2,P3,P4,
  P5,P6,P7,READY,START) );
input CLK,START,B0,B1,B2,B3,A0,A1,A2,A3;
output P4,P5,P6,P7,P0,P1,P2,P3,CNTVCON2,CNTVCO2,READY;

  wire CT2,CNTVG3VD,CT1,CNTVG2VD,CT0,CNTVG1VD,ACVQN3,ACVG4VD1,ACVQN2,ACVG3VD1,ACVQN1,ACVG2VD1,ACVQN0,ACVG1VD1,MRVQN3,MRVG4VD,MRVQN2,MRVG3VD,MRVQN1,MRVG2VD,MRVQN0,MRVG1VD,AX3,AM3,AX2,AM2,AX1,AM1,AX0,AM0,CNTVG3VQN,CNTVG2VQN,CNTVG1VQN,CNTVCON0,CT1N,ACVPCN,CNTVCO0,AMVS0N,IINIIT,READYN,BMVS0N,AMVG5VS0P,AMVG4VS0P,AMVG3VS0P,AMVG2VS0P,AD0,AD0N,AD1,AD1N,AD2,AD2N,AD3,AD3N,CNTVG3VD1,CNTVCON1,CNTVG1VD1,BMVG5VS0P,BMVG4VS0P,BMVG3VS0P,BMVG2VS0P,SMVS0N,ADSH,MRVSHLDN,ADDVC1,ADDVG1VCN,SMVG5VS0P,SMVG4VS0P,SMVG3VS0P,SMVG2VS0P,CNTVG1VZ,CNTVG1VZ1,AMVG5VX,AMVG4VX,AMVG3VX,AMVG2VX,S0,ADDVG1VP,BM3,BMVG5VX,BM2,BMVG4VX,BM1,BMVG3VX,BM0,BMVG2VX,ADDVC2,ADDVG2VCN,S1,ADDVG2VSN,ADDVC3,ADDVG3VCN,S2,ADDVG3VSN,SM0,SMVG2VX,CO,ADDVG4VCN,S3,ADDVG4VSN,SM1,SMVG3VX,SM3,SMVG5VX,SM2,SMVG4VX,AMVG5VG1VAD1NF,AMVG4VG1VAD1NF,AMVG3VG1VAD1NF,AMVG2VG1VAD1NF,BMVG5VG1VAD1NF,BMVG4VG1VAD1NF,BMVG3VG1VAD1NF,BMVG2VG1VAD1NF,AMVG5VG1VAD2NF,AMVG4VG1VAD2NF,AMVG3VG1VAD2NF,AMVG2VG1VAD2NF,ADDVG2VCNVAD1NF,ADDVG3VCNVAD1NF,ADDVG4VCNVAD1NF,MRVG3VDVAD1NF,MRVG2VDVAD1NF,MRVG1VDVAD1NF,BMVG5VG1VAD2NF,BMVG4VG1VAD2NF,BMVG3VG1VAD2NF,BMVG2VG1VAD2NF,SMVG5VG1VAD1NF,SMVG4VG1VAD1NF,SMVG3VG1VAD1NF,SMVG2VG1VAD1NF,ADDVG2VCNVAD4NF,ADDVG2VCNVAD2NF,ADDVG2VCNVOR1NF,MRVG4VDVAD1NF,MRVG4VDVAD2NF,MRVG3VDVAD2NF,MRVG2VDVAD2NF,MRVG1VDVAD2NF,ADDVG2VCNVAD3NF,ADDVG2VCNVOR2NF,ADDVG3VCNVAD4NF,ADDVG3VCNVAD2NF,ADDVG3VCNVOR1NF,ADDVG3VCNVAD3NF,ADDVG3VCNVOR2NF,SMVG2VG1VAD2NF,ADDVG4VCNVAD4NF,ADDVG4VCNVAD2NF,ADDVG4VCNVOR1NF,ADDVG4VCNVAD3NF,ADDVG4VCNVOR2NF,SMVG3VG1VAD2NF,SMVG5VG1VAD2NF,SMVG4VG1VAD2NF,ADDVG1VPVOR1NF,CNTVG3VG2VOR1NF,CNTVG2VG2VOR1NF,CNTVG2VD1,CNTVCO1,CNTVG3VZ1,CNTVG2VZ1,CNTVG3VZ,CNTVG2VZ;

  HS65_LH_DFPRQX4 DFF_0  (.D(CNTVG3VD), .CP(CLK), .RN(a), .Q(CT2) );
  HS65_LH_DFPRQX4 DFF_1 (.D(CNTVG2VD), .CP(CLK), .RN(a), .Q(CT1) );
  HS65_LH_DFPRQX4 DFF_2 (.D(CNTVG1VD), .CP(CLK), .RN(a), .Q(CT0) );
  HS65_LH_DFPRQX4 DFF_3 (.D(ACVG4VD1), .CP(CLK), .RN(a), .Q(ACVQN3) );
  HS65_LH_DFPRQX4 DFF_4 (.D(ACVG3VD1), .CP(CLK), .RN(a), .Q(ACVQN2) );
  HS65_LH_DFPRQX4 DFF_5 (.D(ACVG2VD1), .CP(CLK), .RN(a), .Q(ACVQN1) );
  HS65_LH_DFPRQX4 DFF_6 (.D(ACVG1VD1), .CP(CLK), .RN(a), .Q(ACVQN0) );
  HS65_LH_DFPRQX4 DFF_7 (.D(MRVG4VD), .CP(CLK), .RN(a), .Q(MRVQN3) );
  HS65_LH_DFPRQX4 DFF_8 (.D(MRVG3VD), .CP(CLK), .RN(a), .Q(MRVQN2) );
  HS65_LH_DFPRQX4 DFF_9 (.D(MRVG2VD), .CP(CLK), .RN(a), .Q(MRVQN1) );
  HS65_LH_DFPRQX4 DFF_10 (.D(MRVG1VD), .CP(CLK), .RN(a), .Q(MRVQN0) );
  HS65_LH_DFPRQX4 DFF_11 (.D(AM3), .CP(CLK), .RN(a), .Q(AX3) );
  HS65_LH_DFPRQX4 DFF_12 (.D(AM2), .CP(CLK), .RN(a), .Q(AX2) );
  HS65_LH_DFPRQX4 DFF_13 (.D(AM1), .CP(CLK), .RN(a), .Q(AX1) );
  HS65_LH_DFPRQX4 DFF_14 (.D(AM0), .CP(CLK), .RN(a), .Q(AX0) );
  HS65_LH_IVX2 NOT_0 (.Z(CNTVG3VQN)), .A(CT2) );
  HS65_LH_IVX2 NOT_1 (.Z(CNTVG2VQN), .A(CT1) );
  HS65_LH_IVX2 NOT_2 (.Z(CNTVG1VQN), .A(CT0) );
  HS65_LH_IVX2 NOT_3 (.Z(P7), .A(ACVQN3) );
  HS65_LH_IVX2 NOT_4 (.Z(P6), .A(ACVQN2) );
  HS65_LH_IVX2 NOT_5 (.Z(P5), .A(ACVQN1) );
  HS65_LH_IVX2 NOT_6 (.Z(P4), .A(ACVQN0) );
  HS65_LH_IVX2 NOT_7 (.Z(P3), .A(MRVQN3) );
  HS65_LH_IVX2 NOT_8 (.Z(P2), .A(MRVQN2) );
  HS65_LH_IVX2 NOT_9 (.Z(P1), .A(MRVQN1) );
  HS65_LH_IVX2 NOT_10 (.Z(P0), .A(MRVQN0) );
  HS65_LH_IVX2 NOT_11 (.Z(CNTVCON0), .A(CT0) );
  HS65_LH_IVX2 NOT_12 (.Z(CT1N), .A(CT1) );
  HS65_LH_IVX2 NOT_13 (.Z(ACVPCN), .A(START) );
  HS65_LH_IVX2 NOT_14 (.Z(CNTVCO0), .A(CNTVG1VQN) );
  HS65_LH_IVX2 NOT_15 (.Z(AMVS0N), .A(IINIIT) );
  HS65_LH_IVX2 NOT_16 (.Z(READY), .A(READYN) );
  HS65_LH_IVX2 NOT_17 (.Z(BMVS0N), .A(READYN) );
  HS65_LH_IVX2 NOT_18 (.Z(AMVG5VS0P), .A(AMVS0N) );
  HS65_LH_IVX2 NOT_19 (.Z(AMVG4VS0P), .A(AMVS0N) );
  HS65_LH_IVX2 NOT_20 (.Z(AMVG3VS0P), .A(AMVS0N) );
  HS65_LH_IVX2 NOT_21 (.Z(AMVG2VS0P), .A(AMVS0N) );
  HS65_LH_IVX2 NOT_22 (.Z(AD0), .A(AD0N) );
  HS65_LH_IVX2 NOT_23 (.Z(AD1), .A(AD1N) );
  HS65_LH_IVX2 NOT_24 (.Z(AD2), .A(AD2N) );
  HS65_LH_IVX2 NOT_25 (.Z(AD3), .A(AD3N) );
  HS65_LH_IVX2 NOT_26 (.Z(CNTVG3VD1), .A(CNTVCON1) );
  HS65_LH_IVX2 NOT_27 (.Z(CNTVG1VD1), .A(READY) );
  HS65_LH_IVX2 NOT_28 (.Z(BMVG5VS0P), .A(BMVS0N) );
  HS65_LH_IVX2 NOT_29 (.Z(BMVG4VS0P), .A(BMVS0N) );
  HS65_LH_IVX2 NOT_30 (.Z(BMVG3VS0P), .A(BMVS0N) );
  HS65_LH_IVX2 NOT_31 (.Z(BMVG2VS0P), .A(BMVS0N) );
  HS65_LH_IVX2 NOT_32 (.Z(SMVS0N), .A(ADSH) );
  HS65_LH_IVX2 NOT_33 (.Z(MRVSHLDN), .A(ADSH) );
  HS65_LH_IVX2 NOT_34 (.Z(ADDVC1), .A(ADDVG1VCN) );
  HS65_LH_IVX2 NOT_35 (.Z(SMVG5VS0P), .A(SMVS0N) );
  HS65_LH_IVX2 NOT_36 (.Z(SMVG4VS0P), .A(SMVS0N) );
  HS65_LH_IVX2 NOT_37 (.Z(SMVG3VS0P), .A(SMVS0N) );
  HS65_LH_IVX2 NOT_38 (.Z(SMVG2VS0P), .A(SMVS0N) );
  HS65_LH_IVX2 NOT_39 (.Z(CNTVG1VZ), .A(CNTVG1VZ1) );
  HS65_LH_IVX2 NOT_40 (.Z(AM3), .A(AMVG5VX) );
  HS65_LH_IVX2 NOT_41 (.Z(AM2), .A(AMVG4VX) );
  HS65_LH_IVX2 NOT_42 (.Z(AM1), .A(AMVG3VX) );
  HS65_LH_IVX2 NOT_43 (.Z(AM0), .A(AMVG2VX) );
  HS65_LH_IVX2 NOT_44 (.Z(S0), .A(ADDVG1VP) );
  HS65_LH_IVX2 NOT_45 (.Z(BM3), .A(BMVG5VX) );
  HS65_LH_IVX2 NOT_46 (.Z(BM2), .A(BMVG4VX) );
  HS65_LH_IVX2 NOT_47 (.Z(BM1), .A(BMVG3VX) );
  HS65_LH_IVX2 NOT_48 (.Z(BM0), .A(BMVG2VX) );
  HS65_LH_IVX2 NOT_49 (.Z(ADDVC2), .A(ADDVG2VCN) );
  HS65_LH_IVX2 NOT_50 (.Z(S1), .A(ADDVG2VSN) );
  HS65_LH_IVX2 NOT_51 (.Z(ADDVC3), .A(ADDVG3VCN) );
  HS65_LH_IVX2 NOT_52 (.Z(S2), .A(ADDVG3VSN) );
  HS65_LH_IVX2 NOT_53 (.Z(SM0), .A(SMVG2VX) );
  HS65_LH_IVX2 NOT_54 (.Z(CO), .A(ADDVG4VCN) );
  HS65_LH_IVX2 NOT_55 (.Z(S3), .A(ADDVG4VSN) );
  HS65_LH_IVX2 NOT_56 (.Z(SM1), .A(SMVG3VX) );
  HS65_LH_IVX2 NOT_57 (.Z(SM3), .A(SMVG5VX) );
  HS65_LH_IVX2 NOT_58 (.Z(SM2), .A(SMVG4VX) );
  HS65_LH_AND2X4 AND2_0 (.Z(AMVG5VG1VAD1NF), .A(AMVS0N), .B(AX3) );
  HS65_LH_AND2X4 AND2_1 (.Z(AMVG4VG1VAD1NF), .A(AMVS0N), .B(AX2) );
  HS65_LH_AND2X4 AND2_2 (.Z(AMVG3VG1VAD1NF), .A(AMVS0N), .B(AX1) );
  HS65_LH_AND2X4 AND2_3 (.Z(AMVG2VG1VAD1NF), .A(AMVS0N), .B(AX0) );
  HS65_LH_AND2X4 AND2_4 (.Z(BMVG5VG1VAD1NF), .A(BMVS0N), .B(P3) );
  HS65_LH_AND2X4 AND2_5 (.Z(BMVG4VG1VAD1NF), .A(BMVS0N), .B(P2) );
  HS65_LH_AND2X4 AND2_6 (.Z(BMVG3VG1VAD1NF), .A(BMVS0N), .B(P1) );
  HS65_LH_AND2X4 AND2_7 (.Z(BMVG2VG1VAD1NF), .A(BMVS0N), .B(P0) );
  HS65_LH_AND2X4 AND2_8 (.Z(AMVG5VG1VAD2NF), .A(AMVG5VS0P), .B(A3) );
  HS65_LH_AND2X4 AND2_9 (.Z(AMVG4VG1VAD2NF), .A(AMVG4VS0P), .B(A2) );
  HS65_LH_AND2X4 AND2_10 (.Z(AMVG3VG1VAD2NF), .A(AMVG3VS0P), .B(A1) );
  HS65_LH_AND2X4 AND2_11 (.Z(AMVG2VG1VAD2NF), .A(AMVG2VS0P), .B(A0) );
  HS65_LH_AND2X4 AND2_12 (.Z(ADDVG2VCNVAD1NF), .A(AD1), .B(P5) );
  HS65_LH_AND2X4 AND2_13 (.Z(ADDVG3VCNVAD1NF), .A(AD2), .B(P6) );
  HS65_LH_AND2X4 AND2_14 (.Z(ADDVG4VCNVAD1NF), .A(AD3), .B(P7) );
  HS65_LH_AND2X4 AND2_15 (.Z(MRVG3VDVAD1NF), .A(ADSH), .B(P3) );
  HS65_LH_AND2X4 AND2_16 (.Z(MRVG2VDVAD1NF), .A(ADSH), .B(P2) );
  HS65_LH_AND2X4 AND2_17 (.Z(MRVG1VDVAD1NF), .A(ADSH), .B(P1) );
  HS65_LH_AND2X4 AND2_18 (.Z(BMVG5VG1VAD2NF), .A(BMVG5VS0P), .B(B3) );
  HS65_LH_AND2X4 AND2_19 (.Z(BMVG4VG1VAD2NF), .A(BMVG4VS0P), .B(B2) );
  HS65_LH_AND2X4 AND2_20 (.Z(BMVG3VG1VAD2NF), .A(BMVG3VS0P), .B(B1) );
  HS65_LH_AND2X4 AND2_21 (.Z(BMVG2VG1VAD2NF), .A(BMVG2VS0P), .B(B0) );
  HS65_LH_AND2X4 AND2_22 (.Z(SMVG5VG1VAD1NF), .A(SMVS0N), .B(P7) );
  HS65_LH_AND2X4 AND2_23 (.Z(SMVG4VG1VAD1NF), .A(SMVS0N), .B(P6) );
  HS65_LH_AND2X4 AND2_24 (.Z(SMVG3VG1VAD1NF), .A(SMVS0N), .B(P5) );
  HS65_LH_AND2X4 AND2_25 (.Z(SMVG2VG1VAD1NF), .A(SMVS0N), .B(P4) );
  HS65_LH_AND3X4 AND3_0 (.Z(ADDVG2VCNVAD4NF), .A(ADDVC1), .B(AD1), .C(P5) );
  HS65_LH_AND2X4 AND2_26 (.Z(ADDVG2VCNVAD2NF), .A(ADDVC1), .B(ADDVG2VCNVOR1NF) );
  HS65_LH_AND2X4 AND2_27 (.Z(MRVG4VDVAD1NF), .A(ADSH), .B(S0) );
  HS65_LH_AND2X4 AND2_28 (.Z(MRVG4VDVAD2NF), .A(MRVSHLDN), .B(BM3) );
  HS65_LH_AND2X4 AND2_29 (.Z(MRVG3VDVAD2NF), .A(MRVSHLDN), .B(BM2) );
  HS65_LH_AND2X4 AND2_30 (.Z(MRVG2VDVAD2NF), .A(MRVSHLDN), .B(BM1) );
  HS65_LH_AND2X4 AND2_31 (.Z(MRVG1VDVAD2NF), .A(MRVSHLDN), .B(BM0) );
  HS65_LH_AND2X4 AND2_32 (.Z(ADDVG2VCNVAD3NF), .A(ADDVG2VCNVOR2NF), .B(ADDVG2VCN) );
  HS65_LH_AND3X4 AND3_1 (.Z(ADDVG3VCNVAD4NF), .A(ADDVC2), .B(AD2), .C(P6) );
  HS65_LH_AND2X4 AND2_33 (.Z(ADDVG3VCNVAD2NF), .A(ADDVC2), .B(ADDVG3VCNVOR1NF) );
  HS65_LH_AND2X4 AND2_34 (.Z(ADDVG3VCNVAD3NF), .A(ADDVG3VCNVOR2NF), .B(ADDVG3VCN) );
  HS65_LH_AND2X4 AND2_35 (.Z(SMVG2VG1VAD2NF), .A(SMVG2VS0P), .B(S1) );
  HS65_LH_AND3X4 AND3_2 (.Z(ADDVG4VCNVAD4NF), .A(ADDVC3), .B(AD3), .C(P7) );
  HS65_LH_AND2X4 AND2_36 (.Z(ADDVG4VCNVAD2NF), .A(ADDVC3), .B(ADDVG4VCNVOR1NF) );
  HS65_LH_AND2X4 AND2_37 (.Z(ADDVG4VCNVAD3NF), .A(ADDVG4VCNVOR2NF), .B(ADDVG4VCN) );
  HS65_LH_AND2X4 AND2_38 (.Z(SMVG3VG1VAD2NF), .A(SMVG3VS0P), .B(S2) );
  HS65_LH_AND2X4 AND2_39 (.Z(SMVG5VG1VAD2NF), .A(SMVG5VS0P), .B(CO) );
  HS65_LH_AND2X4 AND2_40 (.Z(SMVG4VG1VAD2NF), .A(SMVG4VS0P), .B(S3) );
  HS65_LH_OR2X4 OR2_0 (.Z(ADDVG1VPVOR1NF), .A(AD0), .B(P4) );
  HS65_LH_OR2X4 OR2_1 (.Z(ADDVG2VCNVOR1NF), .A(AD1), .B(P5) );
  HS65_LH_OR2X4 OR2_2 (.Z(ADDVG3VCNVOR1NF), .A(AD2), .B(P6) );
  HS65_LH_OR2X4 OR2_3 (.Z(ADDVG4VCNVOR1NF), .A(AD3), .B(P7) );
  HS65_LH_OR2X4 OR2_4 (.Z(CNTVG3VG2VOR1NF), .A(CT2), .B(CNTVG3VD1) );
  HS65_LH_OR2X4 OR2_5 (.Z(CNTVG2VG2VOR1NF), .A(CT1), .B(CNTVG2VD1) );
  HS65_LH_OR3X4 OR3_0 (.Z(ADDVG2VCNVOR2NF), .A(ADDVC1), .B(AD1), .C(P5) );
  HS65_LH_OR3X4 OR3_1 (.Z(ADDVG3VCNVOR2NF), .A(ADDVC2), .B(AD2), .C(P6) );
  HS65_LH_OR3X4 OR3_2 (.Z(ADDVG4VCNVOR2NF), .A(ADDVC3), .B(AD3), .C(P7) );
  HS65_LH_NAND3X2 NAND3_0 (.Z(READYN), .A(CT0), .B(CT1N), .C(CT2) );
  HS65_LH_NAND2X2 NAND2_0 (.Z(AD0N), .A(P0), .B(AX0) );
  HS65_LH_NAND2X2 NAND2_1 (.Z(AD1N), .A(P0), .B(AX1) );
  HS65_LH_NAND2X2 NAND2_2 (.Z(AD2N), .A(P0), .B(AX2) );
  HS65_LH_NAND2X2 NAND2_3 (.Z(AD3N), .A(P0), .B(AX3) );
  HS65_LH_NAND2X2 NAND2_4 (.Z(CNTVCON1), .A(CT1), .B(CNTVCO0) );
  HS65_LH_NAND2X2 NAND2_5 (.Z(CNTVCON2), .A(CT2), .B(CNTVCO1) );
  HS65_LH_NAND2X2 NAND2_6 (.Z(ADDVG1VCN), .A(AD0), .B(P4) );
  HS65_LH_NAND2X2 NAND2_7 (.Z(CNTVG3VZ1), .A(CT2), .B(CNTVG3VD1) );
  HS65_LH_NAND2X2 NAND2_8 (.Z(CNTVG2VZ1), .A(CT1), .B(CNTVG2VD1) );
  HS65_LH_NAND2X2 NAND2_9 (.Z(CNTVG1VZ1), .A(CT0), .B(CNTVG1VD1) );
  HS65_LH_NAND2X2 NAND2_10 (.Z(ADDVG1VP), .A(ADDVG1VPVOR1NF), .B(ADDVG1VCN) );
  HS65_LH_NAND2X2 NAND2_11 (.Z(CNTVG3VZ), .A(CNTVG3VG2VOR1NF), .B(CNTVG3VZ1) );
  HS65_LH_NAND2X2 NAND2_12 (.Z(CNTVG2VZ), .A(CNTVG2VG2VOR1NF), .B(CNTVG2VZ1) );
  HS65_LH_NAND2X2 NAND2_13 (.Z(ACVG1VD1), .A(ACVPCN), .B(SM0) );
  HS65_LH_NAND2X2 NAND2_14 (.Z(ACVG2VD1), .A(ACVPCN), .B(SM1) );
  HS65_LH_NAND2X2 NAND2_15 (.Z(ACVG4VD1), .A(ACVPCN), .B(SM3) );
  HS65_LH_NAND2X2 NAND2_16 (.Z(ACVG3VD1), .A(ACVPCN), .B(SM2) );
  HS65_LH_NOR3X2 NOR3_0 (.Z(IINIIT), .A(CT0), .B(CT1), .C(CT2) );
  HS65_LH_NOR2X2 NOR2_0 (.Z(CNTVCO1), .A(CNTVG2VQN), .B(CNTVCON0) );
  HS65_LH_NOR2X2 NOR2_1 (.Z(CNTVCO2), .A(CNTVG3VQN), .B(CNTVCON1) );
  HS65_LH_NOR2X2 NOR2_2 (.Z(ADSH), .A(READY), .B(IINIIT) );
  HS65_LH_NOR2X2 NOR2_3 (.Z(CNTVG2VD1), .A(READY), .B(CNTVCON0) );
  HS65_LH_NOR2X2 NOR2_4 (.Z(AMVG5VX), .A(AMVG5VG1VAD2NF), .B(AMVG5VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_5 (.Z(AMVG4VX), .A(AMVG4VG1VAD2NF), .B(AMVG4VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_6 (.Z(AMVG3VX), .A(AMVG3VG1VAD2NF), .B(AMVG3VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_7 (.Z(AMVG2VX), .A(AMVG2VG1VAD2NF), .B(AMVG2VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_8 (.Z(BMVG5VX), .A(BMVG5VG1VAD2NF), .B(BMVG5VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_9 (.Z(BMVG4VX), .A(BMVG4VG1VAD2NF), .B(BMVG4VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_10 (.Z(BMVG3VX), .A(BMVG3VG1VAD2NF), .B(BMVG3VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_11 (.Z(BMVG2VX), .A(BMVG2VG1VAD2NF), .B(BMVG2VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_12 (.Z(CNTVG3VD), .A(CNTVG3VZ), .B(START) );
  HS65_LH_NOR2X2 NOR2_13 (.Z(CNTVG2VD), .A(CNTVG2VZ), .B(START) );
  HS65_LH_NOR2X2 NOR2_14 (.Z(CNTVG1VD), .A(CNTVG1VZ), .B(START) );
  HS65_LH_NOR2X2 NOR2_15 (.Z(ADDVG2VCN), .A(ADDVG2VCNVAD2NF), .B(ADDVG2VCNVAD1NF) );
  HS65_LH_NOR2X2 NOR2_16 (.Z(MRVG4VD), .A(MRVG4VDVAD2NF), .B(MRVG4VDVAD1NF) );
  HS65_LH_NOR2X2 NOR2_17 (.Z(MRVG3VD), .A(MRVG3VDVAD2NF), .B(MRVG3VDVAD1NF) );
  HS65_LH_NOR2X2 NOR2_18 (.Z(MRVG2VD), .A(MRVG2VDVAD2NF), .B(MRVG2VDVAD1NF) );
  HS65_LH_NOR2X2 NOR2_19 (.Z(MRVG1VD), .A(MRVG1VDVAD2NF), .B(MRVG1VDVAD1NF) );
  HS65_LH_NOR2X2 NOR2_20 (.Z(ADDVG2VSN), .A(ADDVG2VCNVAD4NF), .B(ADDVG2VCNVAD3NF) );
  HS65_LH_NOR2X2 NOR2_21 (.Z(ADDVG3VCN), .A(ADDVG3VCNVAD2NF), .B(ADDVG3VCNVAD1NF) );
  HS65_LH_NOR2X2 NOR2_22 (.Z(ADDVG3VSN), .A(ADDVG3VCNVAD4NF), .B(ADDVG3VCNVAD3NF) );
  HS65_LH_NOR2X2 NOR2_23 (.Z(SMVG2VX), .A(SMVG2VG1VAD2NF), .B(SMVG2VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_24 (.Z(ADDVG4VCN), .A(ADDVG4VCNVAD2NF), .B(ADDVG4VCNVAD1NF) );
  HS65_LH_NOR2X2 NOR2_25 (.Z(ADDVG4VSN), .A(ADDVG4VCNVAD4NF), .B(ADDVG4VCNVAD3NF) );
  HS65_LH_NOR2X2 NOR2_26 (.Z(SMVG3VX), .A(SMVG3VG1VAD2NF), .B(SMVG3VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_27 (.Z(SMVG5VX), .A(SMVG5VG1VAD2NF), .B(SMVG5VG1VAD1NF) );
  HS65_LH_NOR2X2 NOR2_28 (.Z(SMVG4VX), .A(SMVG4VG1VAD2NF), .B(SMVG4VG1VAD1NF) );

endmodule
