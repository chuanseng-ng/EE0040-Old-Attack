module s27(G0,G3);
input G0;
output G3;

  HS65_LH_IVX2 AND2_0 (.Z(G3), .A(G0) );
